-- --------------------------------------------------------------------------------
-- Company : Rochester Institute of Technology (RIT )
-- Engineer : Rohan Patil (rnp5285@rit.edu)
--
-- Create Date : 2/19/19
-- Design Name : instr_mem
-- Module Name : instr_mem - behavioral
-- Project Name : ex3
-- Target Devices : Basys3
--
-- Description :  memory module which holds all instructions to fetch  
-- --------------------------------------------------------------------------------

library IEEE ;
use IEEE . STD_LOGIC_1164 .ALL ;
use IEEE . STD_LOGIC_UNSIGNED .ALL;
use IEEE . NUMERIC_STD .ALL;

entity instr_mem is
    port (
            addr : in std_logic_vector(27 downto 0);
            dout : out std_logic_vector(31 downto 0)
    );
end instr_mem;

architecture behav of instr_mem is
    type mem_type is array(0 to 1023) of std_logic_vector(31 downto 0); -- 2^10 size array, checking the first 10 bits of addr
    -- arbitrary memory values
    signal mem : mem_type := (
        --setup, i type add
        0 => "00100000001000010000000000000010",    -- add r1,r1,#2 = 2
        4 => "00100000010000100000000000000001",    -- add r2,r2,#1 = 1
         -- no op
        8 => "00100000000000000000000000000000",
        12 => "00100000000000000000000000000000",
        16 => "00100000000000000000000000000000",
        20 => "00100000000000000000000000000000",
        -- r type
        -- r1 = 2, r2 = 1
        24 => "00100000010000100000000000000001", -- add r2,r2,#1 = 2
        --24 => "00000000001000100001100000100000", --add r1 + r2 => r3 (3)
        28 => "00000000001000100001100000100100", --and r1 & r2 => r3 (0)
        32 => "00000000001000100001100000011001", --multu r1 * r2 => r3 (2)
        36 => "00000000001000100001100000100101", --or r1 or r2 => r3 (3)
        40 => "00000000001000100001100001000000", --sll r1 sll 1 => r3 (4)
        44 => "00000000001000100001100001000011", --sra r1 sra 1 => r3 (1)
        48 => "00000000001000100001100001000010", --srl r1 srl 1 => r3 (1)
        52 => "00000000001000100001100000100011", --sub r1 - r2 => r3 (1)
        56 => "00000000001000110001100000100000", --add r1 + r3 => r3 (2)
        --56 => "00000000001000100001100000100110", --xor r1 xor r2 => r3 (3)
        -- j type
        60 => "00111100001000010000000000000010", 
        64 => "10001100001000010000000000000010", 
        68 => "00001000000000000000000001000000", -- jump to 256
        256 => "00001100000000000000000000000110", -- jump to 24
        
        --4 => "00100000000000000000000000000000",
--        8 => "00100000000000000000000000000000",
--        12 => "00100000000000000000000000000000",
--        16 => "00100000000000000000000000000000",
--        20 => "00000000001000100001000000100000", --r2 + r1 <= r2
--        24 => "00100000000000000000000000000000",
--        28 => "00100000000000000000000000000000",
--        32 => "00100000000000000000000000000000",
--        36 => "00100000000000000000000000000000",
--        48 => "00000000001000100000100000100000", --r2 + r1 <= r1
--        52 => "00100000000000000000000000000000",
--        56 => "00100000000000000000000000000000",
--        60 => "00100000000000000000000000000000",
--        64 => "00100000000000000000000000000000",
--        68 => "00001000000000000000000000000001", --jump to 4
--        --no-op
--        4 => "00100000000000000000000000000000",
--        8 => "00100000000000000000000000000000",
--        12 => "00100000000000000000000000000000",
--        16 => "00100000000000000000000000000000",
         
        others=>x"00000000"); -- initialize memory location array
begin
    dout <= mem(to_integer(unsigned(addr(9 downto 0))));    -- dout assigned addr idx of mem
end behav;